module ROM(Fatores, Produto);

input [9:0] Fatores;
output [9:0] Produto;

wire [1023:0][9:0] ROM;

assign Produto = ROM[Fatores];

assign 	ROM[{5'd0, 5'd0}] = 10'd0,
	 	ROM[{5'd0, 5'd1}] = 10'd0,
	 	ROM[{5'd0, 5'd2}] = 10'd0,
	 	ROM[{5'd0, 5'd3}] = 10'd0,
	 	ROM[{5'd0, 5'd4}] = 10'd0,
	 	ROM[{5'd0, 5'd5}] = 10'd0,
	 	ROM[{5'd0, 5'd6}] = 10'd0,
	 	ROM[{5'd0, 5'd7}] = 10'd0,
	 	ROM[{5'd0, 5'd8}] = 10'd0,
	 	ROM[{5'd0, 5'd9}] = 10'd0,
	 	ROM[{5'd0, 5'd10}] = 10'd0,
	 	ROM[{5'd0, 5'd11}] = 10'd0,
	 	ROM[{5'd0, 5'd12}] = 10'd0,
	 	ROM[{5'd0, 5'd13}] = 10'd0,
	 	ROM[{5'd0, 5'd14}] = 10'd0,
	 	ROM[{5'd0, 5'd15}] = 10'd0,
	 	ROM[{5'd0, 5'd16}] = 10'd0,
	 	ROM[{5'd0, 5'd17}] = 10'd0,
	 	ROM[{5'd0, 5'd18}] = 10'd0,
	 	ROM[{5'd0, 5'd19}] = 10'd0,
	 	ROM[{5'd0, 5'd20}] = 10'd0,
	 	ROM[{5'd0, 5'd21}] = 10'd0,
	 	ROM[{5'd0, 5'd22}] = 10'd0,
	 	ROM[{5'd0, 5'd23}] = 10'd0,
	 	ROM[{5'd0, 5'd24}] = 10'd0,
	 	ROM[{5'd0, 5'd25}] = 10'd0,
	 	ROM[{5'd0, 5'd26}] = 10'd0,
	 	ROM[{5'd0, 5'd27}] = 10'd0,
	 	ROM[{5'd0, 5'd28}] = 10'd0,
	 	ROM[{5'd0, 5'd29}] = 10'd0,
	 	ROM[{5'd0, 5'd30}] = 10'd0,
	 	ROM[{5'd0, 5'd31}] = 10'd0,
	 	ROM[{5'd1, 5'd0}] = 10'd0,
	 	ROM[{5'd1, 5'd1}] = 10'd1,
	 	ROM[{5'd1, 5'd2}] = 10'd2,
	 	ROM[{5'd1, 5'd3}] = 10'd3,
	 	ROM[{5'd1, 5'd4}] = 10'd4,
	 	ROM[{5'd1, 5'd5}] = 10'd5,
	 	ROM[{5'd1, 5'd6}] = 10'd6,
	 	ROM[{5'd1, 5'd7}] = 10'd7,
	 	ROM[{5'd1, 5'd8}] = 10'd8,
	 	ROM[{5'd1, 5'd9}] = 10'd9,
	 	ROM[{5'd1, 5'd10}] = 10'd10,
	 	ROM[{5'd1, 5'd11}] = 10'd11,
	 	ROM[{5'd1, 5'd12}] = 10'd12,
	 	ROM[{5'd1, 5'd13}] = 10'd13,
	 	ROM[{5'd1, 5'd14}] = 10'd14,
	 	ROM[{5'd1, 5'd15}] = 10'd15,
	 	ROM[{5'd1, 5'd16}] = 10'd16,
	 	ROM[{5'd1, 5'd17}] = 10'd17,
	 	ROM[{5'd1, 5'd18}] = 10'd18,
	 	ROM[{5'd1, 5'd19}] = 10'd19,
	 	ROM[{5'd1, 5'd20}] = 10'd20,
	 	ROM[{5'd1, 5'd21}] = 10'd21,
	 	ROM[{5'd1, 5'd22}] = 10'd22,
	 	ROM[{5'd1, 5'd23}] = 10'd23,
	 	ROM[{5'd1, 5'd24}] = 10'd24,
	 	ROM[{5'd1, 5'd25}] = 10'd25,
	 	ROM[{5'd1, 5'd26}] = 10'd26,
	 	ROM[{5'd1, 5'd27}] = 10'd27,
	 	ROM[{5'd1, 5'd28}] = 10'd28,
	 	ROM[{5'd1, 5'd29}] = 10'd29,
	 	ROM[{5'd1, 5'd30}] = 10'd30,
	 	ROM[{5'd1, 5'd31}] = 10'd31,
	 	ROM[{5'd2, 5'd0}] = 10'd0,
	 	ROM[{5'd2, 5'd1}] = 10'd2,
	 	ROM[{5'd2, 5'd2}] = 10'd4,
	 	ROM[{5'd2, 5'd3}] = 10'd6,
	 	ROM[{5'd2, 5'd4}] = 10'd8,
	 	ROM[{5'd2, 5'd5}] = 10'd10,
	 	ROM[{5'd2, 5'd6}] = 10'd12,
	 	ROM[{5'd2, 5'd7}] = 10'd14,
	 	ROM[{5'd2, 5'd8}] = 10'd16,
	 	ROM[{5'd2, 5'd9}] = 10'd18,
	 	ROM[{5'd2, 5'd10}] = 10'd20,
	 	ROM[{5'd2, 5'd11}] = 10'd22,
	 	ROM[{5'd2, 5'd12}] = 10'd24,
	 	ROM[{5'd2, 5'd13}] = 10'd26,
	 	ROM[{5'd2, 5'd14}] = 10'd28,
	 	ROM[{5'd2, 5'd15}] = 10'd30,
	 	ROM[{5'd2, 5'd16}] = 10'd32,
	 	ROM[{5'd2, 5'd17}] = 10'd34,
	 	ROM[{5'd2, 5'd18}] = 10'd36,
	 	ROM[{5'd2, 5'd19}] = 10'd38,
	 	ROM[{5'd2, 5'd20}] = 10'd40,
	 	ROM[{5'd2, 5'd21}] = 10'd42,
	 	ROM[{5'd2, 5'd22}] = 10'd44,
	 	ROM[{5'd2, 5'd23}] = 10'd46,
	 	ROM[{5'd2, 5'd24}] = 10'd48,
	 	ROM[{5'd2, 5'd25}] = 10'd50,
	 	ROM[{5'd2, 5'd26}] = 10'd52,
	 	ROM[{5'd2, 5'd27}] = 10'd54,
	 	ROM[{5'd2, 5'd28}] = 10'd56,
	 	ROM[{5'd2, 5'd29}] = 10'd58,
	 	ROM[{5'd2, 5'd30}] = 10'd60,
	 	ROM[{5'd2, 5'd31}] = 10'd62,
	 	ROM[{5'd3, 5'd0}] = 10'd0,
	 	ROM[{5'd3, 5'd1}] = 10'd3,
	 	ROM[{5'd3, 5'd2}] = 10'd6,
	 	ROM[{5'd3, 5'd3}] = 10'd9,
	 	ROM[{5'd3, 5'd4}] = 10'd12,
	 	ROM[{5'd3, 5'd5}] = 10'd15,
	 	ROM[{5'd3, 5'd6}] = 10'd18,
	 	ROM[{5'd3, 5'd7}] = 10'd21,
	 	ROM[{5'd3, 5'd8}] = 10'd24,
	 	ROM[{5'd3, 5'd9}] = 10'd27,
	 	ROM[{5'd3, 5'd10}] = 10'd30,
	 	ROM[{5'd3, 5'd11}] = 10'd33,
	 	ROM[{5'd3, 5'd12}] = 10'd36,
	 	ROM[{5'd3, 5'd13}] = 10'd39,
	 	ROM[{5'd3, 5'd14}] = 10'd42,
	 	ROM[{5'd3, 5'd15}] = 10'd45,
	 	ROM[{5'd3, 5'd16}] = 10'd48,
	 	ROM[{5'd3, 5'd17}] = 10'd51,
	 	ROM[{5'd3, 5'd18}] = 10'd54,
	 	ROM[{5'd3, 5'd19}] = 10'd57,
	 	ROM[{5'd3, 5'd20}] = 10'd60,
	 	ROM[{5'd3, 5'd21}] = 10'd63,
	 	ROM[{5'd3, 5'd22}] = 10'd66,
	 	ROM[{5'd3, 5'd23}] = 10'd69,
	 	ROM[{5'd3, 5'd24}] = 10'd72,
	 	ROM[{5'd3, 5'd25}] = 10'd75,
	 	ROM[{5'd3, 5'd26}] = 10'd78,
	 	ROM[{5'd3, 5'd27}] = 10'd81,
	 	ROM[{5'd3, 5'd28}] = 10'd84,
	 	ROM[{5'd3, 5'd29}] = 10'd87,
	 	ROM[{5'd3, 5'd30}] = 10'd90,
	 	ROM[{5'd3, 5'd31}] = 10'd93,
	 	ROM[{5'd4, 5'd0}] = 10'd0,
	 	ROM[{5'd4, 5'd1}] = 10'd4,
	 	ROM[{5'd4, 5'd2}] = 10'd8,
	 	ROM[{5'd4, 5'd3}] = 10'd12,
	 	ROM[{5'd4, 5'd4}] = 10'd16,
	 	ROM[{5'd4, 5'd5}] = 10'd20,
	 	ROM[{5'd4, 5'd6}] = 10'd24,
	 	ROM[{5'd4, 5'd7}] = 10'd28,
	 	ROM[{5'd4, 5'd8}] = 10'd32,
	 	ROM[{5'd4, 5'd9}] = 10'd36,
	 	ROM[{5'd4, 5'd10}] = 10'd40,
	 	ROM[{5'd4, 5'd11}] = 10'd44,
	 	ROM[{5'd4, 5'd12}] = 10'd48,
	 	ROM[{5'd4, 5'd13}] = 10'd52,
	 	ROM[{5'd4, 5'd14}] = 10'd56,
	 	ROM[{5'd4, 5'd15}] = 10'd60,
	 	ROM[{5'd4, 5'd16}] = 10'd64,
	 	ROM[{5'd4, 5'd17}] = 10'd68,
	 	ROM[{5'd4, 5'd18}] = 10'd72,
	 	ROM[{5'd4, 5'd19}] = 10'd76,
	 	ROM[{5'd4, 5'd20}] = 10'd80,
	 	ROM[{5'd4, 5'd21}] = 10'd84,
	 	ROM[{5'd4, 5'd22}] = 10'd88,
	 	ROM[{5'd4, 5'd23}] = 10'd92,
	 	ROM[{5'd4, 5'd24}] = 10'd96,
	 	ROM[{5'd4, 5'd25}] = 10'd100,
	 	ROM[{5'd4, 5'd26}] = 10'd104,
	 	ROM[{5'd4, 5'd27}] = 10'd108,
	 	ROM[{5'd4, 5'd28}] = 10'd112,
	 	ROM[{5'd4, 5'd29}] = 10'd116,
	 	ROM[{5'd4, 5'd30}] = 10'd120,
	 	ROM[{5'd4, 5'd31}] = 10'd124,
	 	ROM[{5'd5, 5'd0}] = 10'd0,
	 	ROM[{5'd5, 5'd1}] = 10'd5,
	 	ROM[{5'd5, 5'd2}] = 10'd10,
	 	ROM[{5'd5, 5'd3}] = 10'd15,
	 	ROM[{5'd5, 5'd4}] = 10'd20,
	 	ROM[{5'd5, 5'd5}] = 10'd25,
	 	ROM[{5'd5, 5'd6}] = 10'd30,
	 	ROM[{5'd5, 5'd7}] = 10'd35,
	 	ROM[{5'd5, 5'd8}] = 10'd40,
	 	ROM[{5'd5, 5'd9}] = 10'd45,
	 	ROM[{5'd5, 5'd10}] = 10'd50,
	 	ROM[{5'd5, 5'd11}] = 10'd55,
	 	ROM[{5'd5, 5'd12}] = 10'd60,
	 	ROM[{5'd5, 5'd13}] = 10'd65,
	 	ROM[{5'd5, 5'd14}] = 10'd70,
	 	ROM[{5'd5, 5'd15}] = 10'd75,
	 	ROM[{5'd5, 5'd16}] = 10'd80,
	 	ROM[{5'd5, 5'd17}] = 10'd85,
	 	ROM[{5'd5, 5'd18}] = 10'd90,
	 	ROM[{5'd5, 5'd19}] = 10'd95,
	 	ROM[{5'd5, 5'd20}] = 10'd100,
	 	ROM[{5'd5, 5'd21}] = 10'd105,
	 	ROM[{5'd5, 5'd22}] = 10'd110,
	 	ROM[{5'd5, 5'd23}] = 10'd115,
	 	ROM[{5'd5, 5'd24}] = 10'd120,
	 	ROM[{5'd5, 5'd25}] = 10'd125,
	 	ROM[{5'd5, 5'd26}] = 10'd130,
	 	ROM[{5'd5, 5'd27}] = 10'd135,
	 	ROM[{5'd5, 5'd28}] = 10'd140,
	 	ROM[{5'd5, 5'd29}] = 10'd145,
	 	ROM[{5'd5, 5'd30}] = 10'd150,
	 	ROM[{5'd5, 5'd31}] = 10'd155,
	 	ROM[{5'd6, 5'd0}] = 10'd0,
	 	ROM[{5'd6, 5'd1}] = 10'd6,
	 	ROM[{5'd6, 5'd2}] = 10'd12,
	 	ROM[{5'd6, 5'd3}] = 10'd18,
	 	ROM[{5'd6, 5'd4}] = 10'd24,
	 	ROM[{5'd6, 5'd5}] = 10'd30,
	 	ROM[{5'd6, 5'd6}] = 10'd36,
	 	ROM[{5'd6, 5'd7}] = 10'd42,
	 	ROM[{5'd6, 5'd8}] = 10'd48,
	 	ROM[{5'd6, 5'd9}] = 10'd54,
	 	ROM[{5'd6, 5'd10}] = 10'd60,
	 	ROM[{5'd6, 5'd11}] = 10'd66,
	 	ROM[{5'd6, 5'd12}] = 10'd72,
	 	ROM[{5'd6, 5'd13}] = 10'd78,
	 	ROM[{5'd6, 5'd14}] = 10'd84,
	 	ROM[{5'd6, 5'd15}] = 10'd90,
	 	ROM[{5'd6, 5'd16}] = 10'd96,
	 	ROM[{5'd6, 5'd17}] = 10'd102,
	 	ROM[{5'd6, 5'd18}] = 10'd108,
	 	ROM[{5'd6, 5'd19}] = 10'd114,
	 	ROM[{5'd6, 5'd20}] = 10'd120,
	 	ROM[{5'd6, 5'd21}] = 10'd126,
	 	ROM[{5'd6, 5'd22}] = 10'd132,
	 	ROM[{5'd6, 5'd23}] = 10'd138,
	 	ROM[{5'd6, 5'd24}] = 10'd144,
	 	ROM[{5'd6, 5'd25}] = 10'd150,
	 	ROM[{5'd6, 5'd26}] = 10'd156,
	 	ROM[{5'd6, 5'd27}] = 10'd162,
	 	ROM[{5'd6, 5'd28}] = 10'd168,
	 	ROM[{5'd6, 5'd29}] = 10'd174,
	 	ROM[{5'd6, 5'd30}] = 10'd180,
	 	ROM[{5'd6, 5'd31}] = 10'd186,
	 	ROM[{5'd7, 5'd0}] = 10'd0,
	 	ROM[{5'd7, 5'd1}] = 10'd7,
	 	ROM[{5'd7, 5'd2}] = 10'd14,
	 	ROM[{5'd7, 5'd3}] = 10'd21,
	 	ROM[{5'd7, 5'd4}] = 10'd28,
	 	ROM[{5'd7, 5'd5}] = 10'd35,
	 	ROM[{5'd7, 5'd6}] = 10'd42,
	 	ROM[{5'd7, 5'd7}] = 10'd49,
	 	ROM[{5'd7, 5'd8}] = 10'd56,
	 	ROM[{5'd7, 5'd9}] = 10'd63,
	 	ROM[{5'd7, 5'd10}] = 10'd70,
	 	ROM[{5'd7, 5'd11}] = 10'd77,
	 	ROM[{5'd7, 5'd12}] = 10'd84,
	 	ROM[{5'd7, 5'd13}] = 10'd91,
	 	ROM[{5'd7, 5'd14}] = 10'd98,
	 	ROM[{5'd7, 5'd15}] = 10'd105,
	 	ROM[{5'd7, 5'd16}] = 10'd112,
	 	ROM[{5'd7, 5'd17}] = 10'd119,
	 	ROM[{5'd7, 5'd18}] = 10'd126,
	 	ROM[{5'd7, 5'd19}] = 10'd133,
	 	ROM[{5'd7, 5'd20}] = 10'd140,
	 	ROM[{5'd7, 5'd21}] = 10'd147,
	 	ROM[{5'd7, 5'd22}] = 10'd154,
	 	ROM[{5'd7, 5'd23}] = 10'd161,
	 	ROM[{5'd7, 5'd24}] = 10'd168,
	 	ROM[{5'd7, 5'd25}] = 10'd175,
	 	ROM[{5'd7, 5'd26}] = 10'd182,
	 	ROM[{5'd7, 5'd27}] = 10'd189,
	 	ROM[{5'd7, 5'd28}] = 10'd196,
	 	ROM[{5'd7, 5'd29}] = 10'd203,
	 	ROM[{5'd7, 5'd30}] = 10'd210,
	 	ROM[{5'd7, 5'd31}] = 10'd217,
	 	ROM[{5'd8, 5'd0}] = 10'd0,
	 	ROM[{5'd8, 5'd1}] = 10'd8,
	 	ROM[{5'd8, 5'd2}] = 10'd16,
	 	ROM[{5'd8, 5'd3}] = 10'd24,
	 	ROM[{5'd8, 5'd4}] = 10'd32,
	 	ROM[{5'd8, 5'd5}] = 10'd40,
	 	ROM[{5'd8, 5'd6}] = 10'd48,
	 	ROM[{5'd8, 5'd7}] = 10'd56,
	 	ROM[{5'd8, 5'd8}] = 10'd64,
	 	ROM[{5'd8, 5'd9}] = 10'd72,
	 	ROM[{5'd8, 5'd10}] = 10'd80,
	 	ROM[{5'd8, 5'd11}] = 10'd88,
	 	ROM[{5'd8, 5'd12}] = 10'd96,
	 	ROM[{5'd8, 5'd13}] = 10'd104,
	 	ROM[{5'd8, 5'd14}] = 10'd112,
	 	ROM[{5'd8, 5'd15}] = 10'd120,
	 	ROM[{5'd8, 5'd16}] = 10'd128,
	 	ROM[{5'd8, 5'd17}] = 10'd136,
	 	ROM[{5'd8, 5'd18}] = 10'd144,
	 	ROM[{5'd8, 5'd19}] = 10'd152,
	 	ROM[{5'd8, 5'd20}] = 10'd160,
	 	ROM[{5'd8, 5'd21}] = 10'd168,
	 	ROM[{5'd8, 5'd22}] = 10'd176,
	 	ROM[{5'd8, 5'd23}] = 10'd184,
	 	ROM[{5'd8, 5'd24}] = 10'd192,
	 	ROM[{5'd8, 5'd25}] = 10'd200,
	 	ROM[{5'd8, 5'd26}] = 10'd208,
	 	ROM[{5'd8, 5'd27}] = 10'd216,
	 	ROM[{5'd8, 5'd28}] = 10'd224,
	 	ROM[{5'd8, 5'd29}] = 10'd232,
	 	ROM[{5'd8, 5'd30}] = 10'd240,
	 	ROM[{5'd8, 5'd31}] = 10'd248,
	 	ROM[{5'd9, 5'd0}] = 10'd0,
	 	ROM[{5'd9, 5'd1}] = 10'd9,
	 	ROM[{5'd9, 5'd2}] = 10'd18,
	 	ROM[{5'd9, 5'd3}] = 10'd27,
	 	ROM[{5'd9, 5'd4}] = 10'd36,
	 	ROM[{5'd9, 5'd5}] = 10'd45,
	 	ROM[{5'd9, 5'd6}] = 10'd54,
	 	ROM[{5'd9, 5'd7}] = 10'd63,
	 	ROM[{5'd9, 5'd8}] = 10'd72,
	 	ROM[{5'd9, 5'd9}] = 10'd81,
	 	ROM[{5'd9, 5'd10}] = 10'd90,
	 	ROM[{5'd9, 5'd11}] = 10'd99,
	 	ROM[{5'd9, 5'd12}] = 10'd108,
	 	ROM[{5'd9, 5'd13}] = 10'd117,
	 	ROM[{5'd9, 5'd14}] = 10'd126,
	 	ROM[{5'd9, 5'd15}] = 10'd135,
	 	ROM[{5'd9, 5'd16}] = 10'd144,
	 	ROM[{5'd9, 5'd17}] = 10'd153,
	 	ROM[{5'd9, 5'd18}] = 10'd162,
	 	ROM[{5'd9, 5'd19}] = 10'd171,
	 	ROM[{5'd9, 5'd20}] = 10'd180,
	 	ROM[{5'd9, 5'd21}] = 10'd189,
	 	ROM[{5'd9, 5'd22}] = 10'd198,
	 	ROM[{5'd9, 5'd23}] = 10'd207,
	 	ROM[{5'd9, 5'd24}] = 10'd216,
	 	ROM[{5'd9, 5'd25}] = 10'd225,
	 	ROM[{5'd9, 5'd26}] = 10'd234,
	 	ROM[{5'd9, 5'd27}] = 10'd243,
	 	ROM[{5'd9, 5'd28}] = 10'd252,
	 	ROM[{5'd9, 5'd29}] = 10'd261,
	 	ROM[{5'd9, 5'd30}] = 10'd270,
	 	ROM[{5'd9, 5'd31}] = 10'd279,
	 	ROM[{5'd10, 5'd0}] = 10'd0,
	 	ROM[{5'd10, 5'd1}] = 10'd10,
	 	ROM[{5'd10, 5'd2}] = 10'd20,
	 	ROM[{5'd10, 5'd3}] = 10'd30,
	 	ROM[{5'd10, 5'd4}] = 10'd40,
	 	ROM[{5'd10, 5'd5}] = 10'd50,
	 	ROM[{5'd10, 5'd6}] = 10'd60,
	 	ROM[{5'd10, 5'd7}] = 10'd70,
	 	ROM[{5'd10, 5'd8}] = 10'd80,
	 	ROM[{5'd10, 5'd9}] = 10'd90,
	 	ROM[{5'd10, 5'd10}] = 10'd100,
	 	ROM[{5'd10, 5'd11}] = 10'd110,
	 	ROM[{5'd10, 5'd12}] = 10'd120,
	 	ROM[{5'd10, 5'd13}] = 10'd130,
	 	ROM[{5'd10, 5'd14}] = 10'd140,
	 	ROM[{5'd10, 5'd15}] = 10'd150,
	 	ROM[{5'd10, 5'd16}] = 10'd160,
	 	ROM[{5'd10, 5'd17}] = 10'd170,
	 	ROM[{5'd10, 5'd18}] = 10'd180,
	 	ROM[{5'd10, 5'd19}] = 10'd190,
	 	ROM[{5'd10, 5'd20}] = 10'd200,
	 	ROM[{5'd10, 5'd21}] = 10'd210,
	 	ROM[{5'd10, 5'd22}] = 10'd220,
	 	ROM[{5'd10, 5'd23}] = 10'd230,
	 	ROM[{5'd10, 5'd24}] = 10'd240,
	 	ROM[{5'd10, 5'd25}] = 10'd250,
	 	ROM[{5'd10, 5'd26}] = 10'd260,
	 	ROM[{5'd10, 5'd27}] = 10'd270,
	 	ROM[{5'd10, 5'd28}] = 10'd280,
	 	ROM[{5'd10, 5'd29}] = 10'd290,
	 	ROM[{5'd10, 5'd30}] = 10'd300,
	 	ROM[{5'd10, 5'd31}] = 10'd310,
	 	ROM[{5'd11, 5'd0}] = 10'd0,
	 	ROM[{5'd11, 5'd1}] = 10'd11,
	 	ROM[{5'd11, 5'd2}] = 10'd22,
	 	ROM[{5'd11, 5'd3}] = 10'd33,
	 	ROM[{5'd11, 5'd4}] = 10'd44,
	 	ROM[{5'd11, 5'd5}] = 10'd55,
	 	ROM[{5'd11, 5'd6}] = 10'd66,
	 	ROM[{5'd11, 5'd7}] = 10'd77,
	 	ROM[{5'd11, 5'd8}] = 10'd88,
	 	ROM[{5'd11, 5'd9}] = 10'd99,
	 	ROM[{5'd11, 5'd10}] = 10'd110,
	 	ROM[{5'd11, 5'd11}] = 10'd121,
	 	ROM[{5'd11, 5'd12}] = 10'd132,
	 	ROM[{5'd11, 5'd13}] = 10'd143,
	 	ROM[{5'd11, 5'd14}] = 10'd154,
	 	ROM[{5'd11, 5'd15}] = 10'd165,
	 	ROM[{5'd11, 5'd16}] = 10'd176,
	 	ROM[{5'd11, 5'd17}] = 10'd187,
	 	ROM[{5'd11, 5'd18}] = 10'd198,
	 	ROM[{5'd11, 5'd19}] = 10'd209,
	 	ROM[{5'd11, 5'd20}] = 10'd220,
	 	ROM[{5'd11, 5'd21}] = 10'd231,
	 	ROM[{5'd11, 5'd22}] = 10'd242,
	 	ROM[{5'd11, 5'd23}] = 10'd253,
	 	ROM[{5'd11, 5'd24}] = 10'd264,
	 	ROM[{5'd11, 5'd25}] = 10'd275,
	 	ROM[{5'd11, 5'd26}] = 10'd286,
	 	ROM[{5'd11, 5'd27}] = 10'd297,
	 	ROM[{5'd11, 5'd28}] = 10'd308,
	 	ROM[{5'd11, 5'd29}] = 10'd319,
	 	ROM[{5'd11, 5'd30}] = 10'd330,
	 	ROM[{5'd11, 5'd31}] = 10'd341,
	 	ROM[{5'd12, 5'd0}] = 10'd0,
	 	ROM[{5'd12, 5'd1}] = 10'd12,
	 	ROM[{5'd12, 5'd2}] = 10'd24,
	 	ROM[{5'd12, 5'd3}] = 10'd36,
	 	ROM[{5'd12, 5'd4}] = 10'd48,
	 	ROM[{5'd12, 5'd5}] = 10'd60,
	 	ROM[{5'd12, 5'd6}] = 10'd72,
	 	ROM[{5'd12, 5'd7}] = 10'd84,
	 	ROM[{5'd12, 5'd8}] = 10'd96,
	 	ROM[{5'd12, 5'd9}] = 10'd108,
	 	ROM[{5'd12, 5'd10}] = 10'd120,
	 	ROM[{5'd12, 5'd11}] = 10'd132,
	 	ROM[{5'd12, 5'd12}] = 10'd144,
	 	ROM[{5'd12, 5'd13}] = 10'd156,
	 	ROM[{5'd12, 5'd14}] = 10'd168,
	 	ROM[{5'd12, 5'd15}] = 10'd180,
	 	ROM[{5'd12, 5'd16}] = 10'd192,
	 	ROM[{5'd12, 5'd17}] = 10'd204,
	 	ROM[{5'd12, 5'd18}] = 10'd216,
	 	ROM[{5'd12, 5'd19}] = 10'd228,
	 	ROM[{5'd12, 5'd20}] = 10'd240,
	 	ROM[{5'd12, 5'd21}] = 10'd252,
	 	ROM[{5'd12, 5'd22}] = 10'd264,
	 	ROM[{5'd12, 5'd23}] = 10'd276,
	 	ROM[{5'd12, 5'd24}] = 10'd288,
	 	ROM[{5'd12, 5'd25}] = 10'd300,
	 	ROM[{5'd12, 5'd26}] = 10'd312,
	 	ROM[{5'd12, 5'd27}] = 10'd324,
	 	ROM[{5'd12, 5'd28}] = 10'd336,
	 	ROM[{5'd12, 5'd29}] = 10'd348,
	 	ROM[{5'd12, 5'd30}] = 10'd360,
	 	ROM[{5'd12, 5'd31}] = 10'd372,
	 	ROM[{5'd13, 5'd0}] = 10'd0,
	 	ROM[{5'd13, 5'd1}] = 10'd13,
	 	ROM[{5'd13, 5'd2}] = 10'd26,
	 	ROM[{5'd13, 5'd3}] = 10'd39,
	 	ROM[{5'd13, 5'd4}] = 10'd52,
	 	ROM[{5'd13, 5'd5}] = 10'd65,
	 	ROM[{5'd13, 5'd6}] = 10'd78,
	 	ROM[{5'd13, 5'd7}] = 10'd91,
	 	ROM[{5'd13, 5'd8}] = 10'd104,
	 	ROM[{5'd13, 5'd9}] = 10'd117,
	 	ROM[{5'd13, 5'd10}] = 10'd130,
	 	ROM[{5'd13, 5'd11}] = 10'd143,
	 	ROM[{5'd13, 5'd12}] = 10'd156,
	 	ROM[{5'd13, 5'd13}] = 10'd169,
	 	ROM[{5'd13, 5'd14}] = 10'd182,
	 	ROM[{5'd13, 5'd15}] = 10'd195,
	 	ROM[{5'd13, 5'd16}] = 10'd208,
	 	ROM[{5'd13, 5'd17}] = 10'd221,
	 	ROM[{5'd13, 5'd18}] = 10'd234,
	 	ROM[{5'd13, 5'd19}] = 10'd247,
	 	ROM[{5'd13, 5'd20}] = 10'd260,
	 	ROM[{5'd13, 5'd21}] = 10'd273,
	 	ROM[{5'd13, 5'd22}] = 10'd286,
	 	ROM[{5'd13, 5'd23}] = 10'd299,
	 	ROM[{5'd13, 5'd24}] = 10'd312,
	 	ROM[{5'd13, 5'd25}] = 10'd325,
	 	ROM[{5'd13, 5'd26}] = 10'd338,
	 	ROM[{5'd13, 5'd27}] = 10'd351,
	 	ROM[{5'd13, 5'd28}] = 10'd364,
	 	ROM[{5'd13, 5'd29}] = 10'd377,
	 	ROM[{5'd13, 5'd30}] = 10'd390,
	 	ROM[{5'd13, 5'd31}] = 10'd403,
	 	ROM[{5'd14, 5'd0}] = 10'd0,
	 	ROM[{5'd14, 5'd1}] = 10'd14,
	 	ROM[{5'd14, 5'd2}] = 10'd28,
	 	ROM[{5'd14, 5'd3}] = 10'd42,
	 	ROM[{5'd14, 5'd4}] = 10'd56,
	 	ROM[{5'd14, 5'd5}] = 10'd70,
	 	ROM[{5'd14, 5'd6}] = 10'd84,
	 	ROM[{5'd14, 5'd7}] = 10'd98,
	 	ROM[{5'd14, 5'd8}] = 10'd112,
	 	ROM[{5'd14, 5'd9}] = 10'd126,
	 	ROM[{5'd14, 5'd10}] = 10'd140,
	 	ROM[{5'd14, 5'd11}] = 10'd154,
	 	ROM[{5'd14, 5'd12}] = 10'd168,
	 	ROM[{5'd14, 5'd13}] = 10'd182,
	 	ROM[{5'd14, 5'd14}] = 10'd196,
	 	ROM[{5'd14, 5'd15}] = 10'd210,
	 	ROM[{5'd14, 5'd16}] = 10'd224,
	 	ROM[{5'd14, 5'd17}] = 10'd238,
	 	ROM[{5'd14, 5'd18}] = 10'd252,
	 	ROM[{5'd14, 5'd19}] = 10'd266,
	 	ROM[{5'd14, 5'd20}] = 10'd280,
	 	ROM[{5'd14, 5'd21}] = 10'd294,
	 	ROM[{5'd14, 5'd22}] = 10'd308,
	 	ROM[{5'd14, 5'd23}] = 10'd322,
	 	ROM[{5'd14, 5'd24}] = 10'd336,
	 	ROM[{5'd14, 5'd25}] = 10'd350,
	 	ROM[{5'd14, 5'd26}] = 10'd364,
	 	ROM[{5'd14, 5'd27}] = 10'd378,
	 	ROM[{5'd14, 5'd28}] = 10'd392,
	 	ROM[{5'd14, 5'd29}] = 10'd406,
	 	ROM[{5'd14, 5'd30}] = 10'd420,
	 	ROM[{5'd14, 5'd31}] = 10'd434,
	 	ROM[{5'd15, 5'd0}] = 10'd0,
	 	ROM[{5'd15, 5'd1}] = 10'd15,
	 	ROM[{5'd15, 5'd2}] = 10'd30,
	 	ROM[{5'd15, 5'd3}] = 10'd45,
	 	ROM[{5'd15, 5'd4}] = 10'd60,
	 	ROM[{5'd15, 5'd5}] = 10'd75,
	 	ROM[{5'd15, 5'd6}] = 10'd90,
	 	ROM[{5'd15, 5'd7}] = 10'd105,
	 	ROM[{5'd15, 5'd8}] = 10'd120,
	 	ROM[{5'd15, 5'd9}] = 10'd135,
	 	ROM[{5'd15, 5'd10}] = 10'd150,
	 	ROM[{5'd15, 5'd11}] = 10'd165,
	 	ROM[{5'd15, 5'd12}] = 10'd180,
	 	ROM[{5'd15, 5'd13}] = 10'd195,
	 	ROM[{5'd15, 5'd14}] = 10'd210,
	 	ROM[{5'd15, 5'd15}] = 10'd225,
	 	ROM[{5'd15, 5'd16}] = 10'd240,
	 	ROM[{5'd15, 5'd17}] = 10'd255,
	 	ROM[{5'd15, 5'd18}] = 10'd270,
	 	ROM[{5'd15, 5'd19}] = 10'd285,
	 	ROM[{5'd15, 5'd20}] = 10'd300,
	 	ROM[{5'd15, 5'd21}] = 10'd315,
	 	ROM[{5'd15, 5'd22}] = 10'd330,
	 	ROM[{5'd15, 5'd23}] = 10'd345,
	 	ROM[{5'd15, 5'd24}] = 10'd360,
	 	ROM[{5'd15, 5'd25}] = 10'd375,
	 	ROM[{5'd15, 5'd26}] = 10'd390,
	 	ROM[{5'd15, 5'd27}] = 10'd405,
	 	ROM[{5'd15, 5'd28}] = 10'd420,
	 	ROM[{5'd15, 5'd29}] = 10'd435,
	 	ROM[{5'd15, 5'd30}] = 10'd450,
	 	ROM[{5'd15, 5'd31}] = 10'd465,
	 	ROM[{5'd16, 5'd0}] = 10'd0,
	 	ROM[{5'd16, 5'd1}] = 10'd16,
	 	ROM[{5'd16, 5'd2}] = 10'd32,
	 	ROM[{5'd16, 5'd3}] = 10'd48,
	 	ROM[{5'd16, 5'd4}] = 10'd64,
	 	ROM[{5'd16, 5'd5}] = 10'd80,
	 	ROM[{5'd16, 5'd6}] = 10'd96,
	 	ROM[{5'd16, 5'd7}] = 10'd112,
	 	ROM[{5'd16, 5'd8}] = 10'd128,
	 	ROM[{5'd16, 5'd9}] = 10'd144,
	 	ROM[{5'd16, 5'd10}] = 10'd160,
	 	ROM[{5'd16, 5'd11}] = 10'd176,
	 	ROM[{5'd16, 5'd12}] = 10'd192,
	 	ROM[{5'd16, 5'd13}] = 10'd208,
	 	ROM[{5'd16, 5'd14}] = 10'd224,
	 	ROM[{5'd16, 5'd15}] = 10'd240,
	 	ROM[{5'd16, 5'd16}] = 10'd256,
	 	ROM[{5'd16, 5'd17}] = 10'd272,
	 	ROM[{5'd16, 5'd18}] = 10'd288,
	 	ROM[{5'd16, 5'd19}] = 10'd304,
	 	ROM[{5'd16, 5'd20}] = 10'd320,
	 	ROM[{5'd16, 5'd21}] = 10'd336,
	 	ROM[{5'd16, 5'd22}] = 10'd352,
	 	ROM[{5'd16, 5'd23}] = 10'd368,
	 	ROM[{5'd16, 5'd24}] = 10'd384,
	 	ROM[{5'd16, 5'd25}] = 10'd400,
	 	ROM[{5'd16, 5'd26}] = 10'd416,
	 	ROM[{5'd16, 5'd27}] = 10'd432,
	 	ROM[{5'd16, 5'd28}] = 10'd448,
	 	ROM[{5'd16, 5'd29}] = 10'd464,
	 	ROM[{5'd16, 5'd30}] = 10'd480,
	 	ROM[{5'd16, 5'd31}] = 10'd496,
	 	ROM[{5'd17, 5'd0}] = 10'd0,
	 	ROM[{5'd17, 5'd1}] = 10'd17,
	 	ROM[{5'd17, 5'd2}] = 10'd34,
	 	ROM[{5'd17, 5'd3}] = 10'd51,
	 	ROM[{5'd17, 5'd4}] = 10'd68,
	 	ROM[{5'd17, 5'd5}] = 10'd85,
	 	ROM[{5'd17, 5'd6}] = 10'd102,
	 	ROM[{5'd17, 5'd7}] = 10'd119,
	 	ROM[{5'd17, 5'd8}] = 10'd136,
	 	ROM[{5'd17, 5'd9}] = 10'd153,
	 	ROM[{5'd17, 5'd10}] = 10'd170,
	 	ROM[{5'd17, 5'd11}] = 10'd187,
	 	ROM[{5'd17, 5'd12}] = 10'd204,
	 	ROM[{5'd17, 5'd13}] = 10'd221,
	 	ROM[{5'd17, 5'd14}] = 10'd238,
	 	ROM[{5'd17, 5'd15}] = 10'd255,
	 	ROM[{5'd17, 5'd16}] = 10'd272,
	 	ROM[{5'd17, 5'd17}] = 10'd289,
	 	ROM[{5'd17, 5'd18}] = 10'd306,
	 	ROM[{5'd17, 5'd19}] = 10'd323,
	 	ROM[{5'd17, 5'd20}] = 10'd340,
	 	ROM[{5'd17, 5'd21}] = 10'd357,
	 	ROM[{5'd17, 5'd22}] = 10'd374,
	 	ROM[{5'd17, 5'd23}] = 10'd391,
	 	ROM[{5'd17, 5'd24}] = 10'd408,
	 	ROM[{5'd17, 5'd25}] = 10'd425,
	 	ROM[{5'd17, 5'd26}] = 10'd442,
	 	ROM[{5'd17, 5'd27}] = 10'd459,
	 	ROM[{5'd17, 5'd28}] = 10'd476,
	 	ROM[{5'd17, 5'd29}] = 10'd493,
	 	ROM[{5'd17, 5'd30}] = 10'd510,
	 	ROM[{5'd17, 5'd31}] = 10'd527,
	 	ROM[{5'd18, 5'd0}] = 10'd0,
	 	ROM[{5'd18, 5'd1}] = 10'd18,
	 	ROM[{5'd18, 5'd2}] = 10'd36,
	 	ROM[{5'd18, 5'd3}] = 10'd54,
	 	ROM[{5'd18, 5'd4}] = 10'd72,
	 	ROM[{5'd18, 5'd5}] = 10'd90,
	 	ROM[{5'd18, 5'd6}] = 10'd108,
	 	ROM[{5'd18, 5'd7}] = 10'd126,
	 	ROM[{5'd18, 5'd8}] = 10'd144,
	 	ROM[{5'd18, 5'd9}] = 10'd162,
	 	ROM[{5'd18, 5'd10}] = 10'd180,
	 	ROM[{5'd18, 5'd11}] = 10'd198,
	 	ROM[{5'd18, 5'd12}] = 10'd216,
	 	ROM[{5'd18, 5'd13}] = 10'd234,
	 	ROM[{5'd18, 5'd14}] = 10'd252,
	 	ROM[{5'd18, 5'd15}] = 10'd270,
	 	ROM[{5'd18, 5'd16}] = 10'd288,
	 	ROM[{5'd18, 5'd17}] = 10'd306,
	 	ROM[{5'd18, 5'd18}] = 10'd324,
	 	ROM[{5'd18, 5'd19}] = 10'd342,
	 	ROM[{5'd18, 5'd20}] = 10'd360,
	 	ROM[{5'd18, 5'd21}] = 10'd378,
	 	ROM[{5'd18, 5'd22}] = 10'd396,
	 	ROM[{5'd18, 5'd23}] = 10'd414,
	 	ROM[{5'd18, 5'd24}] = 10'd432,
	 	ROM[{5'd18, 5'd25}] = 10'd450,
	 	ROM[{5'd18, 5'd26}] = 10'd468,
	 	ROM[{5'd18, 5'd27}] = 10'd486,
	 	ROM[{5'd18, 5'd28}] = 10'd504,
	 	ROM[{5'd18, 5'd29}] = 10'd522,
	 	ROM[{5'd18, 5'd30}] = 10'd540,
	 	ROM[{5'd18, 5'd31}] = 10'd558,
	 	ROM[{5'd19, 5'd0}] = 10'd0,
	 	ROM[{5'd19, 5'd1}] = 10'd19,
	 	ROM[{5'd19, 5'd2}] = 10'd38,
	 	ROM[{5'd19, 5'd3}] = 10'd57,
	 	ROM[{5'd19, 5'd4}] = 10'd76,
	 	ROM[{5'd19, 5'd5}] = 10'd95,
	 	ROM[{5'd19, 5'd6}] = 10'd114,
	 	ROM[{5'd19, 5'd7}] = 10'd133,
	 	ROM[{5'd19, 5'd8}] = 10'd152,
	 	ROM[{5'd19, 5'd9}] = 10'd171,
	 	ROM[{5'd19, 5'd10}] = 10'd190,
	 	ROM[{5'd19, 5'd11}] = 10'd209,
	 	ROM[{5'd19, 5'd12}] = 10'd228,
	 	ROM[{5'd19, 5'd13}] = 10'd247,
	 	ROM[{5'd19, 5'd14}] = 10'd266,
	 	ROM[{5'd19, 5'd15}] = 10'd285,
	 	ROM[{5'd19, 5'd16}] = 10'd304,
	 	ROM[{5'd19, 5'd17}] = 10'd323,
	 	ROM[{5'd19, 5'd18}] = 10'd342,
	 	ROM[{5'd19, 5'd19}] = 10'd361,
	 	ROM[{5'd19, 5'd20}] = 10'd380,
	 	ROM[{5'd19, 5'd21}] = 10'd399,
	 	ROM[{5'd19, 5'd22}] = 10'd418,
	 	ROM[{5'd19, 5'd23}] = 10'd437,
	 	ROM[{5'd19, 5'd24}] = 10'd456,
	 	ROM[{5'd19, 5'd25}] = 10'd475,
	 	ROM[{5'd19, 5'd26}] = 10'd494,
	 	ROM[{5'd19, 5'd27}] = 10'd513,
	 	ROM[{5'd19, 5'd28}] = 10'd532,
	 	ROM[{5'd19, 5'd29}] = 10'd551,
	 	ROM[{5'd19, 5'd30}] = 10'd570,
	 	ROM[{5'd19, 5'd31}] = 10'd589,
	 	ROM[{5'd20, 5'd0}] = 10'd0,
	 	ROM[{5'd20, 5'd1}] = 10'd20,
	 	ROM[{5'd20, 5'd2}] = 10'd40,
	 	ROM[{5'd20, 5'd3}] = 10'd60,
	 	ROM[{5'd20, 5'd4}] = 10'd80,
	 	ROM[{5'd20, 5'd5}] = 10'd100,
	 	ROM[{5'd20, 5'd6}] = 10'd120,
	 	ROM[{5'd20, 5'd7}] = 10'd140,
	 	ROM[{5'd20, 5'd8}] = 10'd160,
	 	ROM[{5'd20, 5'd9}] = 10'd180,
	 	ROM[{5'd20, 5'd10}] = 10'd200,
	 	ROM[{5'd20, 5'd11}] = 10'd220,
	 	ROM[{5'd20, 5'd12}] = 10'd240,
	 	ROM[{5'd20, 5'd13}] = 10'd260,
	 	ROM[{5'd20, 5'd14}] = 10'd280,
	 	ROM[{5'd20, 5'd15}] = 10'd300,
	 	ROM[{5'd20, 5'd16}] = 10'd320,
	 	ROM[{5'd20, 5'd17}] = 10'd340,
	 	ROM[{5'd20, 5'd18}] = 10'd360,
	 	ROM[{5'd20, 5'd19}] = 10'd380,
	 	ROM[{5'd20, 5'd20}] = 10'd400,
	 	ROM[{5'd20, 5'd21}] = 10'd420,
	 	ROM[{5'd20, 5'd22}] = 10'd440,
	 	ROM[{5'd20, 5'd23}] = 10'd460,
	 	ROM[{5'd20, 5'd24}] = 10'd480,
	 	ROM[{5'd20, 5'd25}] = 10'd500,
	 	ROM[{5'd20, 5'd26}] = 10'd520,
	 	ROM[{5'd20, 5'd27}] = 10'd540,
	 	ROM[{5'd20, 5'd28}] = 10'd560,
	 	ROM[{5'd20, 5'd29}] = 10'd580,
	 	ROM[{5'd20, 5'd30}] = 10'd600,
	 	ROM[{5'd20, 5'd31}] = 10'd620,
	 	ROM[{5'd21, 5'd0}] = 10'd0,
	 	ROM[{5'd21, 5'd1}] = 10'd21,
	 	ROM[{5'd21, 5'd2}] = 10'd42,
	 	ROM[{5'd21, 5'd3}] = 10'd63,
	 	ROM[{5'd21, 5'd4}] = 10'd84,
	 	ROM[{5'd21, 5'd5}] = 10'd105,
	 	ROM[{5'd21, 5'd6}] = 10'd126,
	 	ROM[{5'd21, 5'd7}] = 10'd147,
	 	ROM[{5'd21, 5'd8}] = 10'd168,
	 	ROM[{5'd21, 5'd9}] = 10'd189,
	 	ROM[{5'd21, 5'd10}] = 10'd210,
	 	ROM[{5'd21, 5'd11}] = 10'd231,
	 	ROM[{5'd21, 5'd12}] = 10'd252,
	 	ROM[{5'd21, 5'd13}] = 10'd273,
	 	ROM[{5'd21, 5'd14}] = 10'd294,
	 	ROM[{5'd21, 5'd15}] = 10'd315,
	 	ROM[{5'd21, 5'd16}] = 10'd336,
	 	ROM[{5'd21, 5'd17}] = 10'd357,
	 	ROM[{5'd21, 5'd18}] = 10'd378,
	 	ROM[{5'd21, 5'd19}] = 10'd399,
	 	ROM[{5'd21, 5'd20}] = 10'd420,
	 	ROM[{5'd21, 5'd21}] = 10'd441,
	 	ROM[{5'd21, 5'd22}] = 10'd462,
	 	ROM[{5'd21, 5'd23}] = 10'd483,
	 	ROM[{5'd21, 5'd24}] = 10'd504,
	 	ROM[{5'd21, 5'd25}] = 10'd525,
	 	ROM[{5'd21, 5'd26}] = 10'd546,
	 	ROM[{5'd21, 5'd27}] = 10'd567,
	 	ROM[{5'd21, 5'd28}] = 10'd588,
	 	ROM[{5'd21, 5'd29}] = 10'd609,
	 	ROM[{5'd21, 5'd30}] = 10'd630,
	 	ROM[{5'd21, 5'd31}] = 10'd651,
	 	ROM[{5'd22, 5'd0}] = 10'd0,
	 	ROM[{5'd22, 5'd1}] = 10'd22,
	 	ROM[{5'd22, 5'd2}] = 10'd44,
	 	ROM[{5'd22, 5'd3}] = 10'd66,
	 	ROM[{5'd22, 5'd4}] = 10'd88,
	 	ROM[{5'd22, 5'd5}] = 10'd110,
	 	ROM[{5'd22, 5'd6}] = 10'd132,
	 	ROM[{5'd22, 5'd7}] = 10'd154,
	 	ROM[{5'd22, 5'd8}] = 10'd176,
	 	ROM[{5'd22, 5'd9}] = 10'd198,
	 	ROM[{5'd22, 5'd10}] = 10'd220,
	 	ROM[{5'd22, 5'd11}] = 10'd242,
	 	ROM[{5'd22, 5'd12}] = 10'd264,
	 	ROM[{5'd22, 5'd13}] = 10'd286,
	 	ROM[{5'd22, 5'd14}] = 10'd308,
	 	ROM[{5'd22, 5'd15}] = 10'd330,
	 	ROM[{5'd22, 5'd16}] = 10'd352,
	 	ROM[{5'd22, 5'd17}] = 10'd374,
	 	ROM[{5'd22, 5'd18}] = 10'd396,
	 	ROM[{5'd22, 5'd19}] = 10'd418,
	 	ROM[{5'd22, 5'd20}] = 10'd440,
	 	ROM[{5'd22, 5'd21}] = 10'd462,
	 	ROM[{5'd22, 5'd22}] = 10'd484,
	 	ROM[{5'd22, 5'd23}] = 10'd506,
	 	ROM[{5'd22, 5'd24}] = 10'd528,
	 	ROM[{5'd22, 5'd25}] = 10'd550,
	 	ROM[{5'd22, 5'd26}] = 10'd572,
	 	ROM[{5'd22, 5'd27}] = 10'd594,
	 	ROM[{5'd22, 5'd28}] = 10'd616,
	 	ROM[{5'd22, 5'd29}] = 10'd638,
	 	ROM[{5'd22, 5'd30}] = 10'd660,
	 	ROM[{5'd22, 5'd31}] = 10'd682,
	 	ROM[{5'd23, 5'd0}] = 10'd0,
	 	ROM[{5'd23, 5'd1}] = 10'd23,
	 	ROM[{5'd23, 5'd2}] = 10'd46,
	 	ROM[{5'd23, 5'd3}] = 10'd69,
	 	ROM[{5'd23, 5'd4}] = 10'd92,
	 	ROM[{5'd23, 5'd5}] = 10'd115,
	 	ROM[{5'd23, 5'd6}] = 10'd138,
	 	ROM[{5'd23, 5'd7}] = 10'd161,
	 	ROM[{5'd23, 5'd8}] = 10'd184,
	 	ROM[{5'd23, 5'd9}] = 10'd207,
	 	ROM[{5'd23, 5'd10}] = 10'd230,
	 	ROM[{5'd23, 5'd11}] = 10'd253,
	 	ROM[{5'd23, 5'd12}] = 10'd276,
	 	ROM[{5'd23, 5'd13}] = 10'd299,
	 	ROM[{5'd23, 5'd14}] = 10'd322,
	 	ROM[{5'd23, 5'd15}] = 10'd345,
	 	ROM[{5'd23, 5'd16}] = 10'd368,
	 	ROM[{5'd23, 5'd17}] = 10'd391,
	 	ROM[{5'd23, 5'd18}] = 10'd414,
	 	ROM[{5'd23, 5'd19}] = 10'd437,
	 	ROM[{5'd23, 5'd20}] = 10'd460,
	 	ROM[{5'd23, 5'd21}] = 10'd483,
	 	ROM[{5'd23, 5'd22}] = 10'd506,
	 	ROM[{5'd23, 5'd23}] = 10'd529,
	 	ROM[{5'd23, 5'd24}] = 10'd552,
	 	ROM[{5'd23, 5'd25}] = 10'd575,
	 	ROM[{5'd23, 5'd26}] = 10'd598,
	 	ROM[{5'd23, 5'd27}] = 10'd621,
	 	ROM[{5'd23, 5'd28}] = 10'd644,
	 	ROM[{5'd23, 5'd29}] = 10'd667,
	 	ROM[{5'd23, 5'd30}] = 10'd690,
	 	ROM[{5'd23, 5'd31}] = 10'd713,
	 	ROM[{5'd24, 5'd0}] = 10'd0,
	 	ROM[{5'd24, 5'd1}] = 10'd24,
	 	ROM[{5'd24, 5'd2}] = 10'd48,
	 	ROM[{5'd24, 5'd3}] = 10'd72,
	 	ROM[{5'd24, 5'd4}] = 10'd96,
	 	ROM[{5'd24, 5'd5}] = 10'd120,
	 	ROM[{5'd24, 5'd6}] = 10'd144,
	 	ROM[{5'd24, 5'd7}] = 10'd168,
	 	ROM[{5'd24, 5'd8}] = 10'd192,
	 	ROM[{5'd24, 5'd9}] = 10'd216,
	 	ROM[{5'd24, 5'd10}] = 10'd240,
	 	ROM[{5'd24, 5'd11}] = 10'd264,
	 	ROM[{5'd24, 5'd12}] = 10'd288,
	 	ROM[{5'd24, 5'd13}] = 10'd312,
	 	ROM[{5'd24, 5'd14}] = 10'd336,
	 	ROM[{5'd24, 5'd15}] = 10'd360,
	 	ROM[{5'd24, 5'd16}] = 10'd384,
	 	ROM[{5'd24, 5'd17}] = 10'd408,
	 	ROM[{5'd24, 5'd18}] = 10'd432,
	 	ROM[{5'd24, 5'd19}] = 10'd456,
	 	ROM[{5'd24, 5'd20}] = 10'd480,
	 	ROM[{5'd24, 5'd21}] = 10'd504,
	 	ROM[{5'd24, 5'd22}] = 10'd528,
	 	ROM[{5'd24, 5'd23}] = 10'd552,
	 	ROM[{5'd24, 5'd24}] = 10'd576,
	 	ROM[{5'd24, 5'd25}] = 10'd600,
	 	ROM[{5'd24, 5'd26}] = 10'd624,
	 	ROM[{5'd24, 5'd27}] = 10'd648,
	 	ROM[{5'd24, 5'd28}] = 10'd672,
	 	ROM[{5'd24, 5'd29}] = 10'd696,
	 	ROM[{5'd24, 5'd30}] = 10'd720,
	 	ROM[{5'd24, 5'd31}] = 10'd744,
	 	ROM[{5'd25, 5'd0}] = 10'd0,
	 	ROM[{5'd25, 5'd1}] = 10'd25,
	 	ROM[{5'd25, 5'd2}] = 10'd50,
	 	ROM[{5'd25, 5'd3}] = 10'd75,
	 	ROM[{5'd25, 5'd4}] = 10'd100,
	 	ROM[{5'd25, 5'd5}] = 10'd125,
	 	ROM[{5'd25, 5'd6}] = 10'd150,
	 	ROM[{5'd25, 5'd7}] = 10'd175,
	 	ROM[{5'd25, 5'd8}] = 10'd200,
	 	ROM[{5'd25, 5'd9}] = 10'd225,
	 	ROM[{5'd25, 5'd10}] = 10'd250,
	 	ROM[{5'd25, 5'd11}] = 10'd275,
	 	ROM[{5'd25, 5'd12}] = 10'd300,
	 	ROM[{5'd25, 5'd13}] = 10'd325,
	 	ROM[{5'd25, 5'd14}] = 10'd350,
	 	ROM[{5'd25, 5'd15}] = 10'd375,
	 	ROM[{5'd25, 5'd16}] = 10'd400,
	 	ROM[{5'd25, 5'd17}] = 10'd425,
	 	ROM[{5'd25, 5'd18}] = 10'd450,
	 	ROM[{5'd25, 5'd19}] = 10'd475,
	 	ROM[{5'd25, 5'd20}] = 10'd500,
	 	ROM[{5'd25, 5'd21}] = 10'd525,
	 	ROM[{5'd25, 5'd22}] = 10'd550,
	 	ROM[{5'd25, 5'd23}] = 10'd575,
	 	ROM[{5'd25, 5'd24}] = 10'd600,
	 	ROM[{5'd25, 5'd25}] = 10'd625,
	 	ROM[{5'd25, 5'd26}] = 10'd650,
	 	ROM[{5'd25, 5'd27}] = 10'd675,
	 	ROM[{5'd25, 5'd28}] = 10'd700,
	 	ROM[{5'd25, 5'd29}] = 10'd725,
	 	ROM[{5'd25, 5'd30}] = 10'd750,
	 	ROM[{5'd25, 5'd31}] = 10'd775,
	 	ROM[{5'd26, 5'd0}] = 10'd0,
	 	ROM[{5'd26, 5'd1}] = 10'd26,
	 	ROM[{5'd26, 5'd2}] = 10'd52,
	 	ROM[{5'd26, 5'd3}] = 10'd78,
	 	ROM[{5'd26, 5'd4}] = 10'd104,
	 	ROM[{5'd26, 5'd5}] = 10'd130,
	 	ROM[{5'd26, 5'd6}] = 10'd156,
	 	ROM[{5'd26, 5'd7}] = 10'd182,
	 	ROM[{5'd26, 5'd8}] = 10'd208,
	 	ROM[{5'd26, 5'd9}] = 10'd234,
	 	ROM[{5'd26, 5'd10}] = 10'd260,
	 	ROM[{5'd26, 5'd11}] = 10'd286,
	 	ROM[{5'd26, 5'd12}] = 10'd312,
	 	ROM[{5'd26, 5'd13}] = 10'd338,
	 	ROM[{5'd26, 5'd14}] = 10'd364,
	 	ROM[{5'd26, 5'd15}] = 10'd390,
	 	ROM[{5'd26, 5'd16}] = 10'd416,
	 	ROM[{5'd26, 5'd17}] = 10'd442,
	 	ROM[{5'd26, 5'd18}] = 10'd468,
	 	ROM[{5'd26, 5'd19}] = 10'd494,
	 	ROM[{5'd26, 5'd20}] = 10'd520,
	 	ROM[{5'd26, 5'd21}] = 10'd546,
	 	ROM[{5'd26, 5'd22}] = 10'd572,
	 	ROM[{5'd26, 5'd23}] = 10'd598,
	 	ROM[{5'd26, 5'd24}] = 10'd624,
	 	ROM[{5'd26, 5'd25}] = 10'd650,
	 	ROM[{5'd26, 5'd26}] = 10'd676,
	 	ROM[{5'd26, 5'd27}] = 10'd702,
	 	ROM[{5'd26, 5'd28}] = 10'd728,
	 	ROM[{5'd26, 5'd29}] = 10'd754,
	 	ROM[{5'd26, 5'd30}] = 10'd780,
	 	ROM[{5'd26, 5'd31}] = 10'd806,
	 	ROM[{5'd27, 5'd0}] = 10'd0,
	 	ROM[{5'd27, 5'd1}] = 10'd27,
	 	ROM[{5'd27, 5'd2}] = 10'd54,
	 	ROM[{5'd27, 5'd3}] = 10'd81,
	 	ROM[{5'd27, 5'd4}] = 10'd108,
	 	ROM[{5'd27, 5'd5}] = 10'd135,
	 	ROM[{5'd27, 5'd6}] = 10'd162,
	 	ROM[{5'd27, 5'd7}] = 10'd189,
	 	ROM[{5'd27, 5'd8}] = 10'd216,
	 	ROM[{5'd27, 5'd9}] = 10'd243,
	 	ROM[{5'd27, 5'd10}] = 10'd270,
	 	ROM[{5'd27, 5'd11}] = 10'd297,
	 	ROM[{5'd27, 5'd12}] = 10'd324,
	 	ROM[{5'd27, 5'd13}] = 10'd351,
	 	ROM[{5'd27, 5'd14}] = 10'd378,
	 	ROM[{5'd27, 5'd15}] = 10'd405,
	 	ROM[{5'd27, 5'd16}] = 10'd432,
	 	ROM[{5'd27, 5'd17}] = 10'd459,
	 	ROM[{5'd27, 5'd18}] = 10'd486,
	 	ROM[{5'd27, 5'd19}] = 10'd513,
	 	ROM[{5'd27, 5'd20}] = 10'd540,
	 	ROM[{5'd27, 5'd21}] = 10'd567,
	 	ROM[{5'd27, 5'd22}] = 10'd594,
	 	ROM[{5'd27, 5'd23}] = 10'd621,
	 	ROM[{5'd27, 5'd24}] = 10'd648,
	 	ROM[{5'd27, 5'd25}] = 10'd675,
	 	ROM[{5'd27, 5'd26}] = 10'd702,
	 	ROM[{5'd27, 5'd27}] = 10'd729,
	 	ROM[{5'd27, 5'd28}] = 10'd756,
	 	ROM[{5'd27, 5'd29}] = 10'd783,
	 	ROM[{5'd27, 5'd30}] = 10'd810,
	 	ROM[{5'd27, 5'd31}] = 10'd837,
	 	ROM[{5'd28, 5'd0}] = 10'd0,
	 	ROM[{5'd28, 5'd1}] = 10'd28,
	 	ROM[{5'd28, 5'd2}] = 10'd56,
	 	ROM[{5'd28, 5'd3}] = 10'd84,
	 	ROM[{5'd28, 5'd4}] = 10'd112,
	 	ROM[{5'd28, 5'd5}] = 10'd140,
	 	ROM[{5'd28, 5'd6}] = 10'd168,
	 	ROM[{5'd28, 5'd7}] = 10'd196,
	 	ROM[{5'd28, 5'd8}] = 10'd224,
	 	ROM[{5'd28, 5'd9}] = 10'd252,
	 	ROM[{5'd28, 5'd10}] = 10'd280,
	 	ROM[{5'd28, 5'd11}] = 10'd308,
	 	ROM[{5'd28, 5'd12}] = 10'd336,
	 	ROM[{5'd28, 5'd13}] = 10'd364,
	 	ROM[{5'd28, 5'd14}] = 10'd392,
	 	ROM[{5'd28, 5'd15}] = 10'd420,
	 	ROM[{5'd28, 5'd16}] = 10'd448,
	 	ROM[{5'd28, 5'd17}] = 10'd476,
	 	ROM[{5'd28, 5'd18}] = 10'd504,
	 	ROM[{5'd28, 5'd19}] = 10'd532,
	 	ROM[{5'd28, 5'd20}] = 10'd560,
	 	ROM[{5'd28, 5'd21}] = 10'd588,
	 	ROM[{5'd28, 5'd22}] = 10'd616,
	 	ROM[{5'd28, 5'd23}] = 10'd644,
	 	ROM[{5'd28, 5'd24}] = 10'd672,
	 	ROM[{5'd28, 5'd25}] = 10'd700,
	 	ROM[{5'd28, 5'd26}] = 10'd728,
	 	ROM[{5'd28, 5'd27}] = 10'd756,
	 	ROM[{5'd28, 5'd28}] = 10'd784,
	 	ROM[{5'd28, 5'd29}] = 10'd812,
	 	ROM[{5'd28, 5'd30}] = 10'd840,
	 	ROM[{5'd28, 5'd31}] = 10'd868,
	 	ROM[{5'd29, 5'd0}] = 10'd0,
	 	ROM[{5'd29, 5'd1}] = 10'd29,
	 	ROM[{5'd29, 5'd2}] = 10'd58,
	 	ROM[{5'd29, 5'd3}] = 10'd87,
	 	ROM[{5'd29, 5'd4}] = 10'd116,
	 	ROM[{5'd29, 5'd5}] = 10'd145,
	 	ROM[{5'd29, 5'd6}] = 10'd174,
	 	ROM[{5'd29, 5'd7}] = 10'd203,
	 	ROM[{5'd29, 5'd8}] = 10'd232,
	 	ROM[{5'd29, 5'd9}] = 10'd261,
	 	ROM[{5'd29, 5'd10}] = 10'd290,
	 	ROM[{5'd29, 5'd11}] = 10'd319,
	 	ROM[{5'd29, 5'd12}] = 10'd348,
	 	ROM[{5'd29, 5'd13}] = 10'd377,
	 	ROM[{5'd29, 5'd14}] = 10'd406,
	 	ROM[{5'd29, 5'd15}] = 10'd435,
	 	ROM[{5'd29, 5'd16}] = 10'd464,
	 	ROM[{5'd29, 5'd17}] = 10'd493,
	 	ROM[{5'd29, 5'd18}] = 10'd522,
	 	ROM[{5'd29, 5'd19}] = 10'd551,
	 	ROM[{5'd29, 5'd20}] = 10'd580,
	 	ROM[{5'd29, 5'd21}] = 10'd609,
	 	ROM[{5'd29, 5'd22}] = 10'd638,
	 	ROM[{5'd29, 5'd23}] = 10'd667,
	 	ROM[{5'd29, 5'd24}] = 10'd696,
	 	ROM[{5'd29, 5'd25}] = 10'd725,
	 	ROM[{5'd29, 5'd26}] = 10'd754,
	 	ROM[{5'd29, 5'd27}] = 10'd783,
	 	ROM[{5'd29, 5'd28}] = 10'd812,
	 	ROM[{5'd29, 5'd29}] = 10'd841,
	 	ROM[{5'd29, 5'd30}] = 10'd870,
	 	ROM[{5'd29, 5'd31}] = 10'd899,
	 	ROM[{5'd30, 5'd0}] = 10'd0,
	 	ROM[{5'd30, 5'd1}] = 10'd30,
	 	ROM[{5'd30, 5'd2}] = 10'd60,
	 	ROM[{5'd30, 5'd3}] = 10'd90,
	 	ROM[{5'd30, 5'd4}] = 10'd120,
	 	ROM[{5'd30, 5'd5}] = 10'd150,
	 	ROM[{5'd30, 5'd6}] = 10'd180,
	 	ROM[{5'd30, 5'd7}] = 10'd210,
	 	ROM[{5'd30, 5'd8}] = 10'd240,
	 	ROM[{5'd30, 5'd9}] = 10'd270,
	 	ROM[{5'd30, 5'd10}] = 10'd300,
	 	ROM[{5'd30, 5'd11}] = 10'd330,
	 	ROM[{5'd30, 5'd12}] = 10'd360,
	 	ROM[{5'd30, 5'd13}] = 10'd390,
	 	ROM[{5'd30, 5'd14}] = 10'd420,
	 	ROM[{5'd30, 5'd15}] = 10'd450,
	 	ROM[{5'd30, 5'd16}] = 10'd480,
	 	ROM[{5'd30, 5'd17}] = 10'd510,
	 	ROM[{5'd30, 5'd18}] = 10'd540,
	 	ROM[{5'd30, 5'd19}] = 10'd570,
	 	ROM[{5'd30, 5'd20}] = 10'd600,
	 	ROM[{5'd30, 5'd21}] = 10'd630,
	 	ROM[{5'd30, 5'd22}] = 10'd660,
	 	ROM[{5'd30, 5'd23}] = 10'd690,
	 	ROM[{5'd30, 5'd24}] = 10'd720,
	 	ROM[{5'd30, 5'd25}] = 10'd750,
	 	ROM[{5'd30, 5'd26}] = 10'd780,
	 	ROM[{5'd30, 5'd27}] = 10'd810,
	 	ROM[{5'd30, 5'd28}] = 10'd840,
	 	ROM[{5'd30, 5'd29}] = 10'd870,
	 	ROM[{5'd30, 5'd30}] = 10'd900,
	 	ROM[{5'd30, 5'd31}] = 10'd930,
	 	ROM[{5'd31, 5'd0}] = 10'd0,
	 	ROM[{5'd31, 5'd1}] = 10'd31,
	 	ROM[{5'd31, 5'd2}] = 10'd62,
	 	ROM[{5'd31, 5'd3}] = 10'd93,
	 	ROM[{5'd31, 5'd4}] = 10'd124,
	 	ROM[{5'd31, 5'd5}] = 10'd155,
	 	ROM[{5'd31, 5'd6}] = 10'd186,
	 	ROM[{5'd31, 5'd7}] = 10'd217,
	 	ROM[{5'd31, 5'd8}] = 10'd248,
	 	ROM[{5'd31, 5'd9}] = 10'd279,
	 	ROM[{5'd31, 5'd10}] = 10'd310,
	 	ROM[{5'd31, 5'd11}] = 10'd341,
	 	ROM[{5'd31, 5'd12}] = 10'd372,
	 	ROM[{5'd31, 5'd13}] = 10'd403,
	 	ROM[{5'd31, 5'd14}] = 10'd434,
	 	ROM[{5'd31, 5'd15}] = 10'd465,
	 	ROM[{5'd31, 5'd16}] = 10'd496,
	 	ROM[{5'd31, 5'd17}] = 10'd527,
	 	ROM[{5'd31, 5'd18}] = 10'd558,
	 	ROM[{5'd31, 5'd19}] = 10'd589,
	 	ROM[{5'd31, 5'd20}] = 10'd620,
	 	ROM[{5'd31, 5'd21}] = 10'd651,
	 	ROM[{5'd31, 5'd22}] = 10'd682,
	 	ROM[{5'd31, 5'd23}] = 10'd713,
	 	ROM[{5'd31, 5'd24}] = 10'd744,
	 	ROM[{5'd31, 5'd25}] = 10'd775,
	 	ROM[{5'd31, 5'd26}] = 10'd806,
	 	ROM[{5'd31, 5'd27}] = 10'd837,
	 	ROM[{5'd31, 5'd28}] = 10'd868,
	 	ROM[{5'd31, 5'd29}] = 10'd899,
	 	ROM[{5'd31, 5'd30}] = 10'd930,
        ROM[{5'd31, 5'd31}] = 10'd961;

endmodule