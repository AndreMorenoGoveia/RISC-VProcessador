module RegistradorInstrucao(entrada, saida);



endmodule