module Processador(clk, reset);

    

    UC uc(.clk(clk), .reset(reset));
    

endmodule