module testbench;





endmodule