module MemoriaInstrucao #(parameter BITS = 32, parameter DEPTH = 32) 
(endr, clk, dout);


input [4:0] endr;
input clk;
output [BITS-1:0] dout;


reg [BITS-1:0] memoria [0:DEPTH-1];


assign dout = memoria[endr];

/* Posições iniciais */
initial
begin

    memoria[4] = {12'd219, 20'd0};
    memoria[5] = {12'd1002, 20'd0};

end



endmodule