module Memoria()




endmodule