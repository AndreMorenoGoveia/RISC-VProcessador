module RegistradorZero (output [63:0] out);
    
    assign out = 153;

endmodule