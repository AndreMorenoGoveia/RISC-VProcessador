module MemoriaInstrucao 
#(
    parameter BITS = 32,
    parameter DEPTH = 2000,
    parameter i_addr_bits = 6
) 
(addr, dout);


input [i_addr_bits-3:0] addr;
input clk;
output [BITS-1:0] dout;


reg [BITS-1:0] memoria [0:DEPTH-1];


assign dout = memoria[addr];

/* Instruções */
initial
begin

    memoria[0] <= 32'b00000000000000000010000010000011;
    memoria[1] <= 32'b00000000100000000010000100000011;
    memoria[2] <= 32'b00000000000000010000001000110011;
    memoria[3] <= 32'b00000010000100100000001001100011;
    memoria[4] <= 32'b00000000000100100000100001100011;
    memoria[5] <= 32'b00000000000000100000101001100011;
    memoria[6] <= 32'b11111111111100100000001000010011;
    memoria[7] <= 32'b11111110000000000000101011100011;
    memoria[8] <= 32'b01000000000100010000000100110011;
    memoria[9] <= 32'b11111110000000000000001011100011;
    memoria[10] <= 32'b01000000001000001000000010110011;
    memoria[11] <= 32'b11111100000000000000111011100011;
    memoria[12] <= 32'b00000000000100000010100000100011;

end



endmodule