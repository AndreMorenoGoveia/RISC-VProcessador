module Memoria();




endmodule